module xor2 (input wire i0, i1, output wire o);
  assign o = i0 ^ i1;
endmodule 